module clock_divider (
    input wire clk,               // Input clock
    input wire reset,             // Reset signal
    input wire enable,            // Enable signal
    input wire [7:0] div_value,   // 8-bit Divider value
    output reg clk_out            // Output clock
);

    reg [7:0] counter;

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            counter <= 0;
            clk_out <= 0;
        end else if (enable) begin
            if (counter >= div_value) begin
                counter <= 0;
                clk_out <= ~clk_out;
            end else begin
                counter <= counter + 1;
            end
        end
    end
endmodule
